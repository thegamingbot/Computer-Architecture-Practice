module cacheMemory #(
    parameter blocks, words, size
) (
    input clk, 
);
    
endmodule
